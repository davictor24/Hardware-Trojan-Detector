library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity golden_chip is
    Port ( CLK : in STD_LOGIC := '0';
			  CLR : in STD_LOGIC := '0';
           Q : inout STD_LOGIC_VECTOR (9 downto 0) := (others => '0'));
end golden_chip;

architecture Behavioral of golden_chip is
begin
    process(CLK, CLR)
    begin
	     if CLR = '1' then
            Q <= (others => '0');
        elsif rising_edge(CLK) then
            Q <= Q + 1; 
        end if; 
    end process; 

end Behavioral;
